module Phase2();

endmodule